`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/15/2025 12:02:53 AM
// Design Name: 
// Module Name: Definitions
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module Definitions(
`ifndef Multiplexer_Definitions
`define Multiplexer_Definitions
`define Bit_width 16
`endif
    );
endmodule

`ifndef MM_DEFINITIONS_VH
`define MM_DEFINITIONS_VH

`define BIT_WIDTH_DEFAULT  16

`endif
